module NOT_GATE(A,Y);
input A;
output Y;
nor(Y,A);
endmodule
