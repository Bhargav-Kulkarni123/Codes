module Demux_tb;

reg [3:0] S;
wire [15:0] Y;

Demux uut (S,Y);

initial begin

S = 4'b0000; #100;
S = 4'b0001; #100;
S = 4'b0010; #100;
S = 4'b0011; #100;
S = 4'b0100; #100;
S = 4'b0101; #100;
S = 4'b0110; #100;
S = 4'b0111; #100;
S = 4'b1000; #100;
S = 4'b1001; #100;
S = 4'b1010; #100;
S = 4'b1011; #100;
S = 4'b1100; #100;
S = 4'b1101; #100;
S = 4'b1110; #100;
S = 4'b1111; #100;


end
endmodule

