module NOT_GATE(A,Y);
input A;
output Y;
assign Y = ~(A);
endmodule;
